// // Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// // Please do not spread this code without permission 
// module sfp_row (clk, acc, div, fifo_ext_rd, sum_in, sum_out, sfp_in, sfp_out, reset);

//   parameter col = 8;
//   parameter bw = 8;
//   parameter bw_psum = 2*bw+4;

//   input  clk, div, acc, fifo_ext_rd, reset;
//   input  [bw_psum+3:0] sum_in;
//   input  [col*bw_psum-1:0] sfp_in;
//   wire  [col*bw_psum-1:0] abs;
//   reg    div_q;
//   output [col*bw_psum-1:0] sfp_out;
//   output [bw_psum+3:0] sum_out;
//   wire [bw_psum+3:0] sum_this_core;
//   wire [bw_psum+3:0] sum_2core;
//   wire signed [bw_psum-1:0] sfp_in_sign0;
//   wire signed [bw_psum-1:0] sfp_in_sign1;
//   wire signed [bw_psum-1:0] sfp_in_sign2;
//   wire signed [bw_psum-1:0] sfp_in_sign3;
//   wire signed [bw_psum-1:0] sfp_in_sign4;
//   wire signed [bw_psum-1:0] sfp_in_sign5;
//   wire signed [bw_psum-1:0] sfp_in_sign6;
//   wire signed [bw_psum-1:0] sfp_in_sign7;


//   reg [bw_psum+3:0] sfp_out_0;
//   reg [bw_psum+3:0] sfp_out_1;
//   reg [bw_psum+3:0] sfp_out_2;
//   reg [bw_psum+3:0] sfp_out_3;
//   reg [bw_psum+3:0] sfp_out_4;
//   reg [bw_psum+3:0] sfp_out_5;
//   reg [bw_psum+3:0] sfp_out_6;
//   reg [bw_psum+3:0] sfp_out_7;

//   reg [bw_psum+3:0] sum_q;
//   reg fifo_wr;

//   assign sfp_in_sign0 =  sfp_in[bw_psum*1-1 : bw_psum*0];
//   assign sfp_in_sign1 =  sfp_in[bw_psum*2-1 : bw_psum*1];
//   assign sfp_in_sign2 =  sfp_in[bw_psum*3-1 : bw_psum*2];
//   assign sfp_in_sign3 =  sfp_in[bw_psum*4-1 : bw_psum*3];
//   assign sfp_in_sign4 =  sfp_in[bw_psum*5-1 : bw_psum*4];
//   assign sfp_in_sign5 =  sfp_in[bw_psum*6-1 : bw_psum*5];
//   assign sfp_in_sign6 =  sfp_in[bw_psum*7-1 : bw_psum*6];
//   assign sfp_in_sign7 =  sfp_in[bw_psum*8-1 : bw_psum*7];


//   assign sfp_out[bw_psum*1-1 : bw_psum*0] = sfp_out_0;
//   assign sfp_out[bw_psum*2-1 : bw_psum*1] = sfp_out_1;
//   assign sfp_out[bw_psum*3-1 : bw_psum*2] = sfp_out_2;
//   assign sfp_out[bw_psum*4-1 : bw_psum*3] = sfp_out_3;
//   assign sfp_out[bw_psum*5-1 : bw_psum*4] = sfp_out_4;
//   assign sfp_out[bw_psum*6-1 : bw_psum*5] = sfp_out_5;
//   assign sfp_out[bw_psum*7-1 : bw_psum*6] = sfp_out_6;
//   assign sfp_out[bw_psum*8-1 : bw_psum*7] = sfp_out_7;


//   assign sum_2core = sum_this_core + sum_in;

//   assign abs[bw_psum*1-1 : bw_psum*0] = (sfp_in[bw_psum*1-1]) ?  (~sfp_in[bw_psum*1-1 : bw_psum*0] + 1)  :  sfp_in[bw_psum*1-1 : bw_psum*0];
//   assign abs[bw_psum*2-1 : bw_psum*1] = (sfp_in[bw_psum*2-1]) ?  (~sfp_in[bw_psum*2-1 : bw_psum*1] + 1)  :  sfp_in[bw_psum*2-1 : bw_psum*1];
//   assign abs[bw_psum*3-1 : bw_psum*2] = (sfp_in[bw_psum*3-1]) ?  (~sfp_in[bw_psum*3-1 : bw_psum*2] + 1)  :  sfp_in[bw_psum*3-1 : bw_psum*2];
//   assign abs[bw_psum*4-1 : bw_psum*3] = (sfp_in[bw_psum*4-1]) ?  (~sfp_in[bw_psum*4-1 : bw_psum*3] + 1)  :  sfp_in[bw_psum*4-1 : bw_psum*3];
//   assign abs[bw_psum*5-1 : bw_psum*4] = (sfp_in[bw_psum*5-1]) ?  (~sfp_in[bw_psum*5-1 : bw_psum*4] + 1)  :  sfp_in[bw_psum*5-1 : bw_psum*4];
//   assign abs[bw_psum*6-1 : bw_psum*5] = (sfp_in[bw_psum*6-1]) ?  (~sfp_in[bw_psum*6-1 : bw_psum*5] + 1)  :  sfp_in[bw_psum*6-1 : bw_psum*5];
//   assign abs[bw_psum*7-1 : bw_psum*6] = (sfp_in[bw_psum*7-1]) ?  (~sfp_in[bw_psum*7-1 : bw_psum*6] + 1)  :  sfp_in[bw_psum*7-1 : bw_psum*6];
//   assign abs[bw_psum*8-1 : bw_psum*7] = (sfp_in[bw_psum*8-1]) ?  (~sfp_in[bw_psum*8-1 : bw_psum*7] + 1)  :  sfp_in[bw_psum*8-1 : bw_psum*7];

//   wire  full;
//   wire  empty; 


//   fifo #( .DEPTH(6'd32)) fifo_inst_int (
//      .r_clk(clk), 
//      .w_clk(clk), 
//      .i_data(sum_q),
//      .o_data(sum_this_core), 
//      .i_read(div_q), 
//      .i_write(fifo_wr), 
//      .rst(reset),
//      .o_full(full),
// 	   .o_empty(empty)
//   );

//   fifo #( .DEPTH(6'd32)) fifo_inst_ext (
//      .r_clk(clk), 
//      .w_clk(clk), 
//      .i_data(sum_q),
//      .o_data(sum_out), 
//      .i_read(fifo_ext_rd), 
//      .i_write(fifo_wr), 
//      .rst(reset)
//   );

//   // always @(*) begin
//   //   if(fifo_wr) $display("sum_q = %x\n", sum_q);
//   //   if(~fifo_wr && div) $display("sum_this_core = %x\n", sum_this_core);
//   // end

//   always @ (posedge clk) begin
//     if (reset) begin
//       fifo_wr <= 0;
//       div_q <= 0;
//     end
//     else begin
//        div_q <= div ;
//        if (acc) begin
      
//          sum_q <= 
//            {4'b0, abs[bw_psum*1-1 : bw_psum*0]} +
//            {4'b0, abs[bw_psum*2-1 : bw_psum*1]} +
//            {4'b0, abs[bw_psum*3-1 : bw_psum*2]} +
//            {4'b0, abs[bw_psum*4-1 : bw_psum*3]} +
//            {4'b0, abs[bw_psum*5-1 : bw_psum*4]} +
//            {4'b0, abs[bw_psum*6-1 : bw_psum*5]} +
//            {4'b0, abs[bw_psum*7-1 : bw_psum*6]} +
//            {4'b0, abs[bw_psum*8-1 : bw_psum*7]} ;
//          fifo_wr <= 1;
//        end
//        else begin
//          fifo_wr <= 0;
   
//          if (div) begin
//            sfp_out_0 <= (sfp_in[bw_psum*1-1 : bw_psum*0] );
//            sfp_out_1 <= (sfp_in[bw_psum*2-1 : bw_psum*1] );
//            sfp_out_2 <= (sfp_in[bw_psum*3-1 : bw_psum*2] );
//            sfp_out_3 <= (sfp_in[bw_psum*4-1 : bw_psum*3] );
//            sfp_out_4 <= (sfp_in[bw_psum*5-1 : bw_psum*4] );
//            sfp_out_5 <= (sfp_in[bw_psum*6-1 : bw_psum*5] );
//            sfp_out_6 <= (sfp_in[bw_psum*7-1 : bw_psum*6] );
//            sfp_out_7 <= (sfp_in[bw_psum*8-1 : bw_psum*7] );
//           //  $display("sfp_out_sign0 = %x\n", (sfp_out_sign0));

//          end
//        end
//    end
//  end


// endmodule

